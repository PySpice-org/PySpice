* /home/gv/fabrice/developpement/PySpice/examples/spice-parser/kicad-spice-example/kicad-spice-example-0.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: jeu. 26 nov. 2015 16:43:57 CET

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0
* 
* Bring in subckts for power, jacks and opamp
.include components.cir

* Sheet Name: /
U1  Net-_J2-Pad1_ Net-_R1-Pad2_ GND VSS VCC OPAMP		
J1  Net-_J1-Pad1_ GND GND JACK_IN		
J2  Net-_J2-Pad1_ Net-_J2-Pad2_ GND JACK_OUT		
R2  Net-_R1-Pad2_ Net-_J2-Pad1_ 50K		
R1  Net-_J1-Pad1_ Net-_R1-Pad2_ 2K		
R3  GND Net-_J2-Pad2_ 2K		
P1  VSS GND VCC PWR_IN		

.op

.tran 0.1m 3m
.plot tran V(7) V(2)

.ac dec 10 1 100K
.plot ac V(7)

.end
