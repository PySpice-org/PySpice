.title Low Pass RC Filter
Vinput in 0 DC 0V AC SIN(0V 10V 1kHz)
R1 in out 1k
C1 out 0 1u
.ac dec 1 1 10k
.save v(in) v(out)
.control
run
* plot v(out)
print v(out)
.endc
.end
