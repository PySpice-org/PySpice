* **************************************************************************************************

.title STM AN1476: LOW-COST POWER SUPPLY FOR HOME APPLIANCES

* **************************************************************************************************

* 1N4148
.include /home/gv/sys/fc14/fabrice/electronic-design-pattern/spice/libraries/diode/standard-rectifier/1N4148.lib

* 1N5919B: 5.6 V, 3.0 W Zener Diode Voltage Regulator
* d1n5919brl
.include /home/gv/sys/fc14/fabrice/electronic-design-pattern/spice/libraries/diode/zener/1N5919B-spice3.lib

* **************************************************************************************************

.param line_peak_voltage=220V
.param freq=50Hz
.param periode={1 / freq}

Vinput1 out in DC 0V SIN(0V {line_peak_voltage} {freq})
Rload out 0 1k
Cload out 0 220uF
xD1 0 1 1N4148
* xDz1 1 out d1n5919brl
xDz1 1 out 1N4148
Cac 1 2 470nF
Rac 2 in 470

* **************************************************************************************************

.op

.param tran_step={periode / 200}
* .tran 200us 2000ms
.tran {tran_step} {periode * 50}

* **************************************************************************************************

.control
run
plot .1*(V(out)-V(in)), V(out), v(out)-v(1), .1*(V(1)-V(2))
.endc

* **************************************************************************************************

.end

* **************************************************************************************************
