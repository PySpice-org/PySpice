.title ADA4077-2case
* ADA4077-2 SPICE DMod model Typical values
* Description: Amplifier
* Generic Desc: 30V, BIP, OP, Low Noise, Low THD, 2X
* Developed by: RM ADSJ
* Revision History: 02/11/2012 - Updated to new header style
* 0.0 (11/2012)
* Copyright 2008, 2012 by Analog Devices
*
* Refer to "README.DOC" file for License Statement.  Use of this
* model indicates your acceptance of the terms and provisions in
* the License Statement.
*
* Node Assignments
*              noninverting input
*                  |   inverting input
*              |   |   positive supply
*              |   |   |   negative supply
*              |   |   |   |   output
*              |   |   |   |   |
*              |   |   |   |   |
.SUBCKT ADA4077-2   1   2   99   50   45
*#ASSOC Category="Op-amps" symbol=opamp
*
*INPUT STAGE
*
Q1   15 7 60 NIX
Q2   6 2 61 NIX
IOS  1 2 1.75E-10
I1  5 50 77e-6
EOS  7  1 POLY(4) (14,98) (73,98) (81,98) (70,98)  10E-6 1 1 1 1
RC1  11 15 2.6E4
RC2  11 6 2.6E4
RE1 60 5 0.896E2
RE2 61 5 0.896E2
C1   15 6 4.25E-13
D1  50 9 DX
V1  5  9 DC 1.8
D10 99 10 DX
V6 10 11 1.3
*
* CMRR
*
ECM   13 98 POLY(2) (1,98) (2,98) 0 7.192E-4 7.192E-4
RCM1  13 14 2.15E2
RCM2  14 98 5.31E-3
CCM1  13 14 1E-6
*
* PSRR
*
EPSY 72 98 POLY(1) (99,50) -1.683 0.056
CPS3 72 73 1E-6
RPS3 72 73 7.9577E+1
RPS4 73 98 6.5915E-4
*
* EXTRA POLE AND ZERO
*
G1 21 98 (6,15) 26E-6
R1 21 98 9.8E4
R2 21 22 9E6
C2 22 98 1.7614E-12
D3 21 99 DX
D4 50 21 DX
*
* VOLTAGE NOISE
*
VN1 80 98 0
RN1 80 98 16.45E-3
HN  81 98 VN1 6
RN2 81 98 1
*
* FLICKER NOISE
*
D5 69 98 DNOISE
VSN 69 98 DC .60551
H1 70 98 VSN 30.85
RN 70 98 1
*
* INTERNAL VOLTAGE REFERENCE
*
EREF 98  0 POLY(2) (99,0) (50,0) 0 .5 .5
GSY  99 50 POLY(1) (99,50) 130E-6 1.7495E-10
*
* GAIN STAGE
*
G2  98 25 (21,98) 1E-6
R5  25 98 9.9E7
CF  45 25 2.69E-12
V4 25 33 5.3
D7 51 33 DX
EVN 51 98 (50,99) 0.5
V3 32 25 5.3
D6 32 97 DX
EVP 97 98 (99,50) 0.5
*
* OUTPUT STAGE
*
Q3   45 41 99 POUT
Q4   45 43 50 NOUT
RB1  40 41 9.25E4
RB2  42 43 9.25E4
EB1  99 40 POLY(1) (98,25) 0.7153  1
EB2  42 50 POLY(1) (25,98) 0.7153  1
*
* MODELS
*
.MODEL NIX NPN (BF=71429,IS=1E-16)
.MODEL POUT PNP (BF=200,VAF=50,BR=70,IS=1E-15,RC=71.25)
.MODEL NOUT NPN (BF=200,VAF=50,BR=22,IS=1E-15,RC=29.2)
.MODEL DX D(IS=1E-16, RS=5, KF=1E-15)
.MODEL DNOISE D(IS=1E-16,RS=0,KF=1.095E-14)
.ENDS ADA4077-2
*$
Iinj 0 probe 0 AC {0.5*prb*(prb+1)}
Vinj probe Ninplp 0 AC {0.5*prb*(prb-1)}
Vprobe probe Noutlp 0
.model 2N2222 NPN(IS=1E-14 VAF=100
+   BF=200 IKF=0.3 XTB=1.5 BR=3
+   CJC=8E-12 CJE=25E-12 TR=100E-9 TF=400E-12
+   ITF=1 VTF=2 XTF=3 RB=10 RC=.3 RE=.2)
XU1 Ninp Ninn Np15 Nm15 Ninplp ADA4077-2
XU2 No Nre Np15 Nm15 Nrep ADA4077-2
R1 Ninnm 0 {r_1}
R2 Ne Ninnm {r_2}
C2 Ne Ninnm {c_2}
VU1offset Ninn Ninnm {v_1offset}
R3 Nin Ninp {r_3}
VU2offset Nre Nrep {v_2offset}
R4 Nrep Ninp {r_4}
C4 Nrep Ninp {c_4}
R5 Ne No {r_o}
Vi Nin 0 {vin} AC {1-prb*prb}
V2p15 Np15 0 15
Vm15 Nm15 0 -15
Q1 Nc Nb Ne 2N2222
R6 Np15 Nc 50
R7 Noutlp Nb 10
D1 Ngl No YELLOW
Vl Ngl 0 0
.model YELLOW D(IS=93.1P RS=42M N=4.61 BV=2 IBV=10U
+ CJO=2.97P VJ=.75 M=.333 TT=4.32U)
.model NPN NPN
.model PNP PNP
.param prb=0
.param vin=2.5
.param r_1=1k
.param r_2=1k
.param r_3=1k
.param r_4=1k
.param r_o=200
.param c_2=20p
.param c_4=20p
.param v_1offset=0
.param v_2offset=0
.end
