*Sheet Name:/OPA_SR
V1  vp GND dc 1.65 ac 0.5
V2  vn GND dc 1.65 ac -0.5
C2  Vout GND 4p
C1  /3 Vout 6.9p
M7  Vout /6 VDD VDD p_33 W=25.9u L=0.9u
M6  Vout /3 GND GND n_33 W=92.04u L=1.4u
M2  /3 vp /1 VDD p_33 W=51.78u L=0.9u
M1  /2 vn /1 VDD p_33 W=51.78u L=0.9u
M4  /3 /2 GND GND n_33 W=46.02u L=1.4u
M3  /2 /2 GND GND n_33 W=46.02u L=1.4u
M5  /1 /6 VDD VDD p_33 W=12.95u L=0.9u
V0  VDD GND 3.3
M8  /6 /6 VDD VDD p_33 W=1.3u L=0.9u
I1  /6 GND 10u

.lib CMOS_035_Spice_Model.lib tt

.end
