.title Voltage Divider
Vinput in 0 DC 10V
R1 in out 9k
R2 out 0 1k
.op
.end

